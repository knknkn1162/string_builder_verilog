`include "testbench.v"
`include "key_in.v"

module key_in_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
