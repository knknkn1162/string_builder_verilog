`include "testbench.v"
`include "hist_indexer.v"

module hist_indexer_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
