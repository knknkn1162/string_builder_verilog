`include "testbench.v"
`include "posedge_detector.v"

module posedge_detector_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
